
module test(
input	wire    sclk,
input	wire 	rst
);

endmodule